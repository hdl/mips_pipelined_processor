library verilog;
use verilog.vl_types.all;
entity mux_2_1_tb is
end mux_2_1_tb;
