library verilog;
use verilog.vl_types.all;
entity sign_extend_tb is
end sign_extend_tb;
