library verilog;
use verilog.vl_types.all;
entity PC_reg_tb is
end PC_reg_tb;
