library verilog;
use verilog.vl_types.all;
entity register_32_bit_tb is
end register_32_bit_tb;
