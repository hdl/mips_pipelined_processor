library verilog;
use verilog.vl_types.all;
entity processor_tb is
end processor_tb;
